`default_nettype none
`timescale 1ns / 1ps

/* This testbench just instantiates the module and makes some convenient wires
   that can be driven / tested by the cocotb test.py.
*/
module tb ();
   
   // Wire up the inputs and outputs:
   reg clk;
   reg rst_n;
   reg ena;
   reg [7:0] ui_in;
   reg [7:0] uio_in;
   wire [7:0] uo_out;
   wire [7:0] uio_out; 
   wire [7:0] uio_oe;

   wire spi_mosi = uo_out[0];
   wire spi_cs_n = uo_out[1];
   wire spi_clk = uo_out[2];
   wire LEDS = uo_out[3];
	wire TXD = uo_out[4];
   wire spi_clk_ram = uo_out[5];
   wire spi_cs_n_ram = uo_out[6];
   wire spi_mosi_ram = uo_out[7];
   
   assign ui_in [0] = spi_miso;
   assign ui_in [1] = spi_miso_ram;
   assign ui_in [3] = RXD;

`ifdef GL_TEST
  wire VPWR = 1'b1;
  wire VGND = 1'b0;
`endif
   

  // Replace tt_um_example with your module name:
  tt_um_femto user_project (
     `ifdef GL_TEST
     .VPWR(VPWR),
     .VGND(VGND),
     `endif

      .ui_in  (ui_in),    // Dedicated inputs
      .uo_out (uo_out),   // Dedicated outputs
      .uio_in (uio_in),   // IOs: Input path
      .uio_out(uio_out),  // IOs: Output path
      .uio_oe (uio_oe),   // IOs: Enable path (active high: 0=input, 1=output)
      .ena    (ena),      // enable - goes high when design is selected
      .clk    (clk),      // clock
      .rst_n  (rst_n)     // not reset
  );

endmodule
